module execute(
	// Inputs
	setDataZero,pc_as_operand,currPC,SrcA,SrcB,alu_op,immValue,immSel,addConstant4,
	//Outputs
	alu_out
	);
///////////////////////////////////////
/////////////// Inputs ///////////////
/////////////////////////////////////
input setDataZero,pc_as_operand,immSel,addConstant4;
input [31:0]currPC,SrcA,SrcB,immValue;
input [4:0] alu_op;
////////////////////////////////////////
/////////////// Outputs ///////////////
//////////////////////////////////////
output [31:0] alu_out;

//////////////////////////////////////////
/////////////// Variables ///////////////
////////////////////////////////////////

logic [31:0] alu_inA,alu_inB;

////////////////////////////////////////
///////////////////////////////////////
//////////////////////////////////////

assign alu_inA = (setDataZero) ? 32'h0 : (pc_as_operand) ? currPC : SrcA;
assign alu_inB = (addConstant4) ? 32'h4 : (immSel) ? immValue : SrcB;




endmodule
