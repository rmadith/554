/*
    CS/ECE 552 Spring '23
    Eric Dubberstein, Joash Shankar

    256 bit decoder
*/
`default_nettype none
module decoder8to256(
    // inputs
    index, enable, 
    
    // output
    decoder_out);

    input wire enable;
    input wire [7:0] index;
    output wire decoder_out;
	
	reg decoder_out_i;
	
	always@(*) begin
		case(index)
			8'd0: decoder_out_i = 256'd1;
			8'd1: decoder_out_i = 256'd2;
			8'd2: decoder_out_i = 256'd4;
			8'd3: decoder_out_i = 256'd8;
			8'd4: decoder_out_i = 256'd16;
			8'd5: decoder_out_i = 256'd32;
			8'd6: decoder_out_i = 256'd64;
			8'd7: decoder_out_i = 256'd128;
			8'd8: decoder_out_i = 256'd256;
			8'd9: decoder_out_i = 256'd512;
			8'd10: decoder_out_i = 256'd1024;
			8'd11: decoder_out_i = 256'd2048;
			8'd12: decoder_out_i = 256'd4096;
			8'd13: decoder_out_i = 256'd8192;
			8'd14: decoder_out_i = 256'd16384;
			8'd15: decoder_out_i = 256'd32768;
			8'd16: decoder_out_i = 256'd65536;
			8'd17: decoder_out_i = 256'd131072;
			8'd18: decoder_out_i = 256'd262144;
			8'd19: decoder_out_i = 256'd524288;
			8'd20: decoder_out_i = 256'd1048576;
			8'd21: decoder_out_i = 256'd2097152;
			8'd22: decoder_out_i = 256'd4194304;
			8'd23: decoder_out_i = 256'd8388608;
			8'd24: decoder_out_i = 256'd16777216;
			8'd25: decoder_out_i = 256'd33554432;
			8'd26: decoder_out_i = 256'd67108864;
			8'd27: decoder_out_i = 256'd134217728;
			8'd28: decoder_out_i = 256'd268435456;
			8'd29: decoder_out_i = 256'd536870912;
			8'd30: decoder_out_i = 256'd1073741824;
			8'd31: decoder_out_i = 256'd2147483648;
			8'd32: decoder_out_i = 256'd4294967296;
			8'd33: decoder_out_i = 256'd8589934592;
			8'd34: decoder_out_i = 256'd17179869184;
			8'd35: decoder_out_i = 256'd34359738368;
			8'd36: decoder_out_i = 256'd68719476736;
			8'd37: decoder_out_i = 256'd137438953472;
			8'd38: decoder_out_i = 256'd274877906944;
			8'd39: decoder_out_i = 256'd549755813888;
			8'd40: decoder_out_i = 256'd1099511627776;
			8'd41: decoder_out_i = 256'd2199023255552;
			8'd42: decoder_out_i = 256'd4398046511104;
			8'd43: decoder_out_i = 256'd8796093022208;
			8'd44: decoder_out_i = 256'd17592186044416;
			8'd45: decoder_out_i = 256'd35184372088832;
			8'd46: decoder_out_i = 256'd70368744177664;
			8'd47: decoder_out_i = 256'd140737488355328;
			8'd48: decoder_out_i = 256'd281474976710656;
			8'd49: decoder_out_i = 256'd562949953421312;
			8'd50: decoder_out_i = 256'd1125899906842624;
			8'd51: decoder_out_i = 256'd2251799813685248;
			8'd52: decoder_out_i = 256'd4503599627370496;
			8'd53: decoder_out_i = 256'd9007199254740992;
			8'd54: decoder_out_i = 256'd18014398509481984;
			8'd55: decoder_out_i = 256'd36028797018963968;
			8'd56: decoder_out_i = 256'd72057594037927936;
			8'd57: decoder_out_i = 256'd144115188075855872;
			8'd58: decoder_out_i = 256'd288230376151711744;
			8'd59: decoder_out_i = 256'd576460752303423488;
			8'd60: decoder_out_i = 256'd1152921504606846976;
			8'd61: decoder_out_i = 256'd2305843009213693952;
			8'd62: decoder_out_i = 256'd4611686018427387904;
			8'd63: decoder_out_i = 256'd9223372036854775808;
			8'd64: decoder_out_i = 256'd18446744073709551616;
			8'd65: decoder_out_i = 256'd36893488147419103232;
			8'd66: decoder_out_i = 256'd73786976294838206464;
			8'd67: decoder_out_i = 256'd147573952589676412928;
			8'd68: decoder_out_i = 256'd295147905179352825856;
			8'd69: decoder_out_i = 256'd590295810358705651712;
			8'd70: decoder_out_i = 256'd1180591620717411303424;
			8'd71: decoder_out_i = 256'd2361183241434822606848;
			8'd72: decoder_out_i = 256'd4722366482869645213696;
			8'd73: decoder_out_i = 256'd9444732965739290427392;
			8'd74: decoder_out_i = 256'd18889465931478580854784;
			8'd75: decoder_out_i = 256'd37778931862957161709568;
			8'd76: decoder_out_i = 256'd75557863725914323419136;
			8'd77: decoder_out_i = 256'd151115727451828646838272;
			8'd78: decoder_out_i = 256'd302231454903657293676544;
			8'd79: decoder_out_i = 256'd604462909807314587353088;
			8'd80: decoder_out_i = 256'd1208925819614629174706176;
			8'd81: decoder_out_i = 256'd2417851639229258349412352;
			8'd82: decoder_out_i = 256'd4835703278458516698824704;
			8'd83: decoder_out_i = 256'd9671406556917033397649408;
			8'd84: decoder_out_i = 256'd19342813113834066795298816;
			8'd85: decoder_out_i = 256'd38685626227668133590597632;
			8'd86: decoder_out_i = 256'd77371252455336267181195264;
			8'd87: decoder_out_i = 256'd154742504910672534362390528;
			8'd88: decoder_out_i = 256'd309485009821345068724781056;
			8'd89: decoder_out_i = 256'd618970019642690137449562112;
			8'd90: decoder_out_i = 256'd1237940039285380274899124224;
			8'd91: decoder_out_i = 256'd2475880078570760549798248448;
			8'd92: decoder_out_i = 256'd4951760157141521099596496896;
			8'd93: decoder_out_i = 256'd9903520314283042199192993792;
			8'd94: decoder_out_i = 256'd19807040628566084398385987584;
			8'd95: decoder_out_i = 256'd39614081257132168796771975168;
			8'd96: decoder_out_i = 256'd79228162514264337593543950336;
			8'd97: decoder_out_i = 256'd158456325028528675187087900672;
			8'd98: decoder_out_i = 256'd316912650057057350374175801344;
			8'd99: decoder_out_i = 256'd633825300114114700748351602688;
			8'd100: decoder_out_i = 256'd1267650600228229401496703205376;
			8'd101: decoder_out_i = 256'd2535301200456458802993406410752;
			8'd102: decoder_out_i = 256'd5070602400912917605986812821504;
			8'd103: decoder_out_i = 256'd10141204801825835211973625643008;
			8'd104: decoder_out_i = 256'd20282409603651670423947251286016;
			8'd105: decoder_out_i = 256'd40564819207303340847894502572032;
			8'd106: decoder_out_i = 256'd81129638414606681695789005144064;
			8'd107: decoder_out_i = 256'd162259276829213363391578010288128;
			8'd108: decoder_out_i = 256'd324518553658426726783156020576256;
			8'd109: decoder_out_i = 256'd649037107316853453566312041152512;
			8'd110: decoder_out_i = 256'd1298074214633706907132624082305024;
			8'd111: decoder_out_i = 256'd2596148429267413814265248164610048;
			8'd112: decoder_out_i = 256'd5192296858534827628530496329220096;
			8'd113: decoder_out_i = 256'd10384593717069655257060992658440192;
			8'd114: decoder_out_i = 256'd20769187434139310514121985316880384;
			8'd115: decoder_out_i = 256'd41538374868278621028243970633760768;
			8'd116: decoder_out_i = 256'd83076749736557242056487941267521536;
			8'd117: decoder_out_i = 256'd166153499473114484112975882535043072;
			8'd118: decoder_out_i = 256'd332306998946228968225951765070086144;
			8'd119: decoder_out_i = 256'd664613997892457936451903530140172288;
			8'd120: decoder_out_i = 256'd1329227995784915872903807060280344576;
			8'd121: decoder_out_i = 256'd2658455991569831745807614120560689152;
			8'd122: decoder_out_i = 256'd5316911983139663491615228241121378304;
			8'd123: decoder_out_i = 256'd10633823966279326983230456482242756608;
			8'd124: decoder_out_i = 256'd21267647932558653966460912964485513216;
			8'd125: decoder_out_i = 256'd42535295865117307932921825928971026432;
			8'd126: decoder_out_i = 256'd85070591730234615865843651857942052864;
			8'd127: decoder_out_i = 256'd170141183460469231731687303715884105728;
			8'd128: decoder_out_i = 256'd340282366920938463463374607431768211456;
			8'd129: decoder_out_i = 256'd680564733841876926926749214863536422912;
			8'd130: decoder_out_i = 256'd1361129467683753853853498429727072845824;
			8'd131: decoder_out_i = 256'd2722258935367507707706996859454145691648;
			8'd132: decoder_out_i = 256'd5444517870735015415413993718908291383296;
			8'd133: decoder_out_i = 256'd10889035741470030830827987437816582766592;
			8'd134: decoder_out_i = 256'd21778071482940061661655974875633165533184;
			8'd135: decoder_out_i = 256'd43556142965880123323311949751266331066368;
			8'd136: decoder_out_i = 256'd87112285931760246646623899502532662132736;
			8'd137: decoder_out_i = 256'd174224571863520493293247799005065324265472;
			8'd138: decoder_out_i = 256'd348449143727040986586495598010130648530944;
			8'd139: decoder_out_i = 256'd696898287454081973172991196020261297061888;
			8'd140: decoder_out_i = 256'd1393796574908163946345982392040522594123776;
			8'd141: decoder_out_i = 256'd2787593149816327892691964784081045188247552;
			8'd142: decoder_out_i = 256'd5575186299632655785383929568162090376495104;
			8'd143: decoder_out_i = 256'd11150372599265311570767859136324180752990208;
			8'd144: decoder_out_i = 256'd22300745198530623141535718272648361505980416;
			8'd145: decoder_out_i = 256'd44601490397061246283071436545296723011960832;
			8'd146: decoder_out_i = 256'd89202980794122492566142873090593446023921664;
			8'd147: decoder_out_i = 256'd178405961588244985132285746181186892047843328;
			8'd148: decoder_out_i = 256'd356811923176489970264571492362373784095686656;
			8'd149: decoder_out_i = 256'd713623846352979940529142984724747568191373312;
			8'd150: decoder_out_i = 256'd1427247692705959881058285969449495136382746624;
			8'd151: decoder_out_i = 256'd2854495385411919762116571938898990272765493248;
			8'd152: decoder_out_i = 256'd5708990770823839524233143877797980545530986496;
			8'd153: decoder_out_i = 256'd11417981541647679048466287755595961091061972992;
			8'd154: decoder_out_i = 256'd22835963083295358096932575511191922182123945984;
			8'd155: decoder_out_i = 256'd45671926166590716193865151022383844364247891968;
			8'd156: decoder_out_i = 256'd91343852333181432387730302044767688728495783936;
			8'd157: decoder_out_i = 256'd182687704666362864775460604089535377456991567872;
			8'd158: decoder_out_i = 256'd365375409332725729550921208179070754913983135744;
			8'd159: decoder_out_i = 256'd730750818665451459101842416358141509827966271488;
			8'd160: decoder_out_i = 256'd1461501637330902918203684832716283019655932542976;
			8'd161: decoder_out_i = 256'd2923003274661805836407369665432566039311865085952;
			8'd162: decoder_out_i = 256'd5846006549323611672814739330865132078623730171904;
			8'd163: decoder_out_i = 256'd11692013098647223345629478661730264157247460343808;
			8'd164: decoder_out_i = 256'd23384026197294446691258957323460528314494920687616;
			8'd165: decoder_out_i = 256'd46768052394588893382517914646921056628989841375232;
			8'd166: decoder_out_i = 256'd93536104789177786765035829293842113257979682750464;
			8'd167: decoder_out_i = 256'd187072209578355573530071658587684226515959365500928;
			8'd168: decoder_out_i = 256'd374144419156711147060143317175368453031918731001856;
			8'd169: decoder_out_i = 256'd748288838313422294120286634350736906063837462003712;
			8'd170: decoder_out_i = 256'd1496577676626844588240573268701473812127674924007424;
			8'd171: decoder_out_i = 256'd2993155353253689176481146537402947624255349848014848;
			8'd172: decoder_out_i = 256'd5986310706507378352962293074805895248510699696029696;
			8'd173: decoder_out_i = 256'd11972621413014756705924586149611790497021399392059392;
			8'd174: decoder_out_i = 256'd23945242826029513411849172299223580994042798784118784;
			8'd175: decoder_out_i = 256'd47890485652059026823698344598447161988085597568237568;
			8'd176: decoder_out_i = 256'd95780971304118053647396689196894323976171195136475136;
			8'd177: decoder_out_i = 256'd191561942608236107294793378393788647952342390272950272;
			8'd178: decoder_out_i = 256'd383123885216472214589586756787577295904684780545900544;
			8'd179: decoder_out_i = 256'd766247770432944429179173513575154591809369561091801088;
			8'd180: decoder_out_i = 256'd1532495540865888858358347027150309183618739122183602176;
			8'd181: decoder_out_i = 256'd3064991081731777716716694054300618367237478244367204352;
			8'd182: decoder_out_i = 256'd6129982163463555433433388108601236734474956488734408704;
			8'd183: decoder_out_i = 256'd12259964326927110866866776217202473468949912977468817408;
			8'd184: decoder_out_i = 256'd24519928653854221733733552434404946937899825954937634816;
			8'd185: decoder_out_i = 256'd49039857307708443467467104868809893875799651909875269632;
			8'd186: decoder_out_i = 256'd98079714615416886934934209737619787751599303819750539264;
			8'd187: decoder_out_i = 256'd196159429230833773869868419475239575503198607639501078528;
			8'd188: decoder_out_i = 256'd392318858461667547739736838950479151006397215279002157056;
			8'd189: decoder_out_i = 256'd784637716923335095479473677900958302012794430558004314112;
			8'd190: decoder_out_i = 256'd1569275433846670190958947355801916604025588861116008628224;
			8'd191: decoder_out_i = 256'd3138550867693340381917894711603833208051177722232017256448;
			8'd192: decoder_out_i = 256'd6277101735386680763835789423207666416102355444464034512896;
			8'd193: decoder_out_i = 256'd12554203470773361527671578846415332832204710888928069025792;
			8'd194: decoder_out_i = 256'd25108406941546723055343157692830665664409421777856138051584;
			8'd195: decoder_out_i = 256'd50216813883093446110686315385661331328818843555712276103168;
			8'd196: decoder_out_i = 256'd100433627766186892221372630771322662657637687111424552206336;
			8'd197: decoder_out_i = 256'd200867255532373784442745261542645325315275374222849104412672;
			8'd198: decoder_out_i = 256'd401734511064747568885490523085290650630550748445698208825344;
			8'd199: decoder_out_i = 256'd803469022129495137770981046170581301261101496891396417650688;
			8'd200: decoder_out_i = 256'd1606938044258990275541962092341162602522202993782792835301376;
			8'd201: decoder_out_i = 256'd3213876088517980551083924184682325205044405987565585670602752;
			8'd202: decoder_out_i = 256'd6427752177035961102167848369364650410088811975131171341205504;
			8'd203: decoder_out_i = 256'd12855504354071922204335696738729300820177623950262342682411008;
			8'd204: decoder_out_i = 256'd25711008708143844408671393477458601640355247900524685364822016;
			8'd205: decoder_out_i = 256'd51422017416287688817342786954917203280710495801049370729644032;
			8'd206: decoder_out_i = 256'd102844034832575377634685573909834406561420991602098741459288064;
			8'd207: decoder_out_i = 256'd205688069665150755269371147819668813122841983204197482918576128;
			8'd208: decoder_out_i = 256'd411376139330301510538742295639337626245683966408394965837152256;
			8'd209: decoder_out_i = 256'd822752278660603021077484591278675252491367932816789931674304512;
			8'd210: decoder_out_i = 256'd1645504557321206042154969182557350504982735865633579863348609024;
			8'd211: decoder_out_i = 256'd3291009114642412084309938365114701009965471731267159726697218048;
			8'd212: decoder_out_i = 256'd6582018229284824168619876730229402019930943462534319453394436096;
			8'd213: decoder_out_i = 256'd13164036458569648337239753460458804039861886925068638906788872192;
			8'd214: decoder_out_i = 256'd26328072917139296674479506920917608079723773850137277813577744384;
			8'd215: decoder_out_i = 256'd52656145834278593348959013841835216159447547700274555627155488768;
			8'd216: decoder_out_i = 256'd105312291668557186697918027683670432318895095400549111254310977536;
			8'd217: decoder_out_i = 256'd210624583337114373395836055367340864637790190801098222508621955072;
			8'd218: decoder_out_i = 256'd421249166674228746791672110734681729275580381602196445017243910144;
			8'd219: decoder_out_i = 256'd842498333348457493583344221469363458551160763204392890034487820288;
			8'd220: decoder_out_i = 256'd1684996666696914987166688442938726917102321526408785780068975640576;
			8'd221: decoder_out_i = 256'd3369993333393829974333376885877453834204643052817571560137951281152;
			8'd222: decoder_out_i = 256'd6739986666787659948666753771754907668409286105635143120275902562304;
			8'd223: decoder_out_i = 256'd13479973333575319897333507543509815336818572211270286240551805124608;
			8'd224: decoder_out_i = 256'd26959946667150639794667015087019630673637144422540572481103610249216;
			8'd225: decoder_out_i = 256'd53919893334301279589334030174039261347274288845081144962207220498432;
			8'd226: decoder_out_i = 256'd107839786668602559178668060348078522694548577690162289924414440996864;
			8'd227: decoder_out_i = 256'd215679573337205118357336120696157045389097155380324579848828881993728;
			8'd228: decoder_out_i = 256'd431359146674410236714672241392314090778194310760649159697657763987456;
			8'd229: decoder_out_i = 256'd862718293348820473429344482784628181556388621521298319395315527974912;
			8'd230: decoder_out_i = 256'd1725436586697640946858688965569256363112777243042596638790631055949824;
			8'd231: decoder_out_i = 256'd3450873173395281893717377931138512726225554486085193277581262111899648;
			8'd232: decoder_out_i = 256'd6901746346790563787434755862277025452451108972170386555162524223799296;
			8'd233: decoder_out_i = 256'd13803492693581127574869511724554050904902217944340773110325048447598592;
			8'd234: decoder_out_i = 256'd27606985387162255149739023449108101809804435888681546220650096895197184;
			8'd235: decoder_out_i = 256'd55213970774324510299478046898216203619608871777363092441300193790394368;
			8'd236: decoder_out_i = 256'd110427941548649020598956093796432407239217743554726184882600387580788736;
			8'd237: decoder_out_i = 256'd220855883097298041197912187592864814478435487109452369765200775161577472;
			8'd238: decoder_out_i = 256'd441711766194596082395824375185729628956870974218904739530401550323154944;
			8'd239: decoder_out_i = 256'd883423532389192164791648750371459257913741948437809479060803100646309888;
			8'd240: decoder_out_i = 256'd1766847064778384329583297500742918515827483896875618958121606201292619776;
			8'd241: decoder_out_i = 256'd3533694129556768659166595001485837031654967793751237916243212402585239552;
			8'd242: decoder_out_i = 256'd7067388259113537318333190002971674063309935587502475832486424805170479104;
			8'd243: decoder_out_i = 256'd14134776518227074636666380005943348126619871175004951664972849610340958208;
			8'd244: decoder_out_i = 256'd28269553036454149273332760011886696253239742350009903329945699220681916416;
			8'd245: decoder_out_i = 256'd56539106072908298546665520023773392506479484700019806659891398441363832832;
			8'd246: decoder_out_i = 256'd113078212145816597093331040047546785012958969400039613319782796882727665664;
			8'd247: decoder_out_i = 256'd226156424291633194186662080095093570025917938800079226639565593765455331328;
			8'd248: decoder_out_i = 256'd452312848583266388373324160190187140051835877600158453279131187530910662656;
			8'd249: decoder_out_i = 256'd904625697166532776746648320380374280103671755200316906558262375061821325312;
			8'd250: decoder_out_i = 256'd1809251394333065553493296640760748560207343510400633813116524750123642650624;
			8'd251: decoder_out_i = 256'd3618502788666131106986593281521497120414687020801267626233049500247285301248;
			8'd252: decoder_out_i = 256'd7237005577332262213973186563042994240829374041602535252466099000494570602496;
			8'd253: decoder_out_i = 256'd14474011154664524427946373126085988481658748083205070504932198000989141204992;
			8'd254: decoder_out_i = 256'd28948022309329048855892746252171976963317496166410141009864396001978282409984;
			8'd255: decoder_out_i = 256'd57896044618658097711785492504343953926634992332820282019728792003956564819968; 
		endcase
	end
	
	assign decoder_out = decoder_out_i & enable;

endmodule
`default_nettype wire
