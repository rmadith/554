`default_nettype none

module cpu(
	input wire logic clk, 
	input wire logic rst_n

);

	/////////////// fetch (outputs) //////////////////
	logic [31:0] PC_plus4_IFID_in;
	logic [31:0] instruction_IFID_in;
    logic [31:0] PC_IFID_in;
	logic ECALL_IFID_in;

	/////////////// IFID pipeline register (outputs) //////////////////
	logic [31:0] PC_plus4_IFID_out;
	logic [31:0] instruction_IFID_IDEX;
    logic [31:0] PC_IFID_IDEX;
	logic ECALL_IFID_IDEX;

	////////////////// decode (outputs) //////////////////
	logic [31:0] regData1_IDEX_in;
	logic [31:0] regData2_IDEX_in;
	logic [31:0] sext_imm_IDEX_in;

	logic immSel_IDEX_in;
	logic PC_as_operand_IDEX_in;
	logic setDataZero_IDEX_in;
	logic [3:0] ALU_op_IDEX_in;
	logic memRead_IDEX_in; 
	logic [2:0] memType_IDEX_in; 
	logic memWrite_IDEX_in;
	logic addConstant4_IDEX_in;
	logic regWriteEnable_IDEX_in;

	logic [31:0] branch_PC;
	logic takeBranch;

	/////////////// IDEX pipeline register (outputs) //////////////////
	logic [31:0] regData1_IDEX_out;
	logic [31:0] regData2_IDEX_out;
	logic [31:0] sext_imm_IDEX_out;

	logic immSel_IDEX_out;
	logic PC_as_operand_IDEX_out;
	logic setDataZero_IDEX_out;
	logic [3:0] ALU_op_IDEX_out;
	logic memRead_IDEX_EXMEM; 
	logic [2:0] memType_IDEX_EXMEM; 
	logic memWrite_IDEX_EXMEM;
	logic addConstant4_IDEX_out;
	logic regWriteEnable_IDEX_EXMEM;

	logic [31:0] instruction_IDEX_EXMEM;
	logic [31:0] PC_IDEX_EXMEM;

	logic ECALL_IDEX_EXMEM;

	////////////////// execute (outputs) //////////////////
	logic [31:0] execute_result_EXMEM_in;


	/////////////// EXMEM pipeline register (outputs) //////////////////
	logic regWriteEnable_EXMEM_MEMWB;
    logic [31:0] instruction_EXMEM_MEMWB;
    logic [31:0] PC_EXMEM_MEMWB;
    logic [31:0] regData2_EXMEM_out;
    logic [2:0] memType_EXMEM_out;
    logic memRead_EXMEM_MEMWB;
    logic memWrite_EXMEM_out;
    logic [31:0] execute_result_EXMEM_MEMWB;
	logic ECALL_EXMEM_MEMWB;


	////////////////// memory (outputs) //////////////////
	logic [31:0] memReadRst_MEMWB_in;

	/////////////// MEMWB pipeline register (outputs) //////////////////
	logic regWriteEnable_MEMWB_out;
    logic [31:0] instruction_MEMWB_out;
    logic [31:0] PC_MEMWB_out;
    logic [31:0] execute_result_MEMWB_out;
    logic memRead_MEMWB_out;
    logic [31:0] memReadRst_MEMWB_out;
	logic ECALL_MEMWB_out;

	////////////////// writeback (outputs) //////////////////
	logic [31:0] writeBackData;



	// Instantiate the modules for each stage of (what will be) the pipeline.
	fetch iFetch(
		///// INPUTS  /////
		.clk(clk),
		.rst_n(rst_n),

		.PC_enable(1'b1), 
		.takeBranch(takeBranch),
		.branch_PC(branch_PC), 
		.incorrect_b_prediction(1'b0),
		.PC_IFID_IDEX(PC_IFID_IDEX),
		.PC_plus4_IFID_out(PC_plus4_IFID_out),

		///// OUTPUTS /////
		.PC_plus4_IFID_in(PC_plus4_IFID_in),
		.instruction_IFID_in(instruction_IFID_in),
		.PC_IFID_in(PC_IFID_in), 
		.ECALL(ECALL_IFID_in)
    );

	IFIDpipelineReg iIFID_pipeline_reg(
		///// INPUTS  /////
		.clk(clk),
		.rst_n(rst_n),
		.stall_disable(1'b0),
		.flush(1'b0),

		///// PIPELINE INPUTS  /////
		.PC_plus4_IFID_in(PC_plus4_IFID_in),
		.instruction_IFID_in(instruction_IFID_in),
		.PC_IFID_in(PC_IFID_in),
		.ECALL_IFID_in(ECALL_IFID_in),

		///// PIPELINE OUTPUTS  /////
		.PC_plus4_IFID_out(PC_plus4_IFID_out),
		.instruction_IFID_IDEX(instruction_IFID_IDEX),
		.PC_IFID_IDEX(PC_IFID_IDEX), 
		.ECALL_IFID_IDEX(ECALL_IFID_IDEX)
	);
	

	decode iDecode(
		///// INPUTS  /////
		.clk(clk),
		.rst_n(rst_n),

		.instruction_IFID_IDEX(instruction_IFID_IDEX),
		.PC_IFID_IDEX(PC_IFID_IDEX),
		.PC_plus4_IFID_out(PC_plus4_IFID_out),

		.instruction_MEMWB_out(instruction_MEMWB_out),
		.writeBackData(writeBackData),
		

		///// OUTPUTS /////
		.regData1_IDEX_in(regData1_IDEX_in),
		.regData2_IDEX_in(regData2_IDEX_in),
		.sext_imm_IDEX_in(sext_imm_IDEX_in),

		.immSel_IDEX_in(immSel_IDEX_in),
		.PC_as_operand_IDEX_in(PC_as_operand_IDEX_in),
		.setDataZero_IDEX_in(setDataZero_IDEX_in),
		.ALU_op_IDEX_in(ALU_op_IDEX_in),
		.memRead_IDEX_in(memRead_IDEX_in),
		.memType_IDEX_in(memType_IDEX_in),
		.memWrite_IDEX_in(memWrite_IDEX_in),
		.addConstant4_IDEX_in(addConstant4_IDEX_in),
		.regWriteEnable_IDEX_in(regWriteEnable_IDEX_in),

		.branch_PC(branch_PC),
		.takeBranch(takeBranch)
	);

	IDEXpipelineReg iIDEX_pipeline_reg(
		///// INPUTS  /////
		.clk(clk),
		.rst_n(rst_n),
		
		.stall_disable(1'b0),
		.flush(1'b0),

		///// PIPELINE INPUTS  /////
		.regData1_IDEX_in(regData1_IDEX_in),
		.regData2_IDEX_in(regData2_IDEX_in),
		.sext_imm_IDEX_in(sext_imm_IDEX_in),

		.immSel_IDEX_in(immSel_IDEX_in),
		.PC_as_operand_IDEX_in(PC_as_operand_IDEX_in),
		.setDataZero_IDEX_in(setDataZero_IDEX_in),
		.ALU_op_IDEX_in(ALU_op_IDEX_in),
		.memRead_IDEX_in(memRead_IDEX_in), 
		.memType_IDEX_in(memType_IDEX_in), 
		.memWrite_IDEX_in(memWrite_IDEX_in),
		.addConstant4_IDEX_in(addConstant4_IDEX_in),
		.regWriteEnable_IDEX_in(regWriteEnable_IDEX_in),

		.instruction_IFID_IDEX(instruction_IFID_IDEX),
		.PC_IFID_IDEX(PC_IFID_IDEX),
		.ECALL_IFID_IDEX(ECALL_IFID_IDEX),


		///// PIPELINE OUTPUTS  /////
		.regData1_IDEX_out(regData1_IDEX_out),
		.regData2_IDEX_out(regData2_IDEX_out),
		.sext_imm_IDEX_out(sext_imm_IDEX_out),

		.immSel_IDEX_out(immSel_IDEX_out),
		.PC_as_operand_IDEX_out(PC_as_operand_IDEX_out),
		.setDataZero_IDEX_out(setDataZero_IDEX_out),
		.ALU_op_IDEX_out(ALU_op_IDEX_out),
		.memRead_IDEX_EXMEM(memRead_IDEX_EXMEM), 
		.memType_IDEX_EXMEM(memType_IDEX_EXMEM), 
		.memWrite_IDEX_EXMEM(memWrite_IDEX_EXMEM),
		.addConstant4_IDEX_out(addConstant4_IDEX_out),
		.regWriteEnable_IDEX_EXMEM(regWriteEnable_IDEX_EXMEM),

		.instruction_IDEX_EXMEM(instruction_IDEX_EXMEM),
		.PC_IDEX_EXMEM(PC_IDEX_EXMEM), 

		.ECALL_IDEX_EXMEM(ECALL_IDEX_EXMEM)

	);

	


	execute iExecute(
		///// INPUTS  /////
		.setDataZero_IDEX_out(setDataZero_IDEX_out),
		.PC_as_operand_IDEX_out(PC_as_operand_IDEX_out),
		.regData1_IDEX_out(regData1_IDEX_out),
		.regData2_IDEX_out(regData2_IDEX_out),
		.immSel_IDEX_out(immSel_IDEX_out),
		.sext_imm_IDEX_out(sext_imm_IDEX_out),
		.ALU_op_IDEX_out(ALU_op_IDEX_out),
		.PC_IDEX_EXMEM(PC_IDEX_EXMEM),
		.memRead_IDEX_EXMEM(memRead_IDEX_EXMEM),
		.memWrite_IDEX_EXMEM(memWrite_IDEX_EXMEM),
		.addConstant4_IDEX_out(addConstant4_IDEX_out),

		///// OUTPUTS  /////
		.execute_result_EXMEM_in(execute_result_EXMEM_in)
	);

	EXMEMpipelineReg iEXMEM_pipeline_reg(
		///// INPUTS  /////
		.clk(clk),
		.rst_n(rst_n),
		
		.stall_disable(1'b0),
		.flush(1'b0),

		///// PIPELINE INPUTS  /////
		.regWriteEnable_IDEX_EXMEM(regWriteEnable_IDEX_EXMEM),
		.instruction_IDEX_EXMEM(instruction_IDEX_EXMEM),
		.PC_IDEX_EXMEM(PC_IDEX_EXMEM),
		.regData2_EXMEM_in(regData2_IDEX_out), // NOTE: will be connected to output of forwarding unit eventually.
		.memType_IDEX_EXMEM(memType_IDEX_EXMEM),
		.memRead_IDEX_EXMEM(memRead_IDEX_EXMEM),
		.memWrite_IDEX_EXMEM(memWrite_IDEX_EXMEM),
		.execute_result_EXMEM_in(execute_result_EXMEM_in),
		.ECALL_IDEX_EXMEM(ECALL_IDEX_EXMEM),

		///// PIPELINE OUTPUTS  /////
		.regWriteEnable_EXMEM_MEMWB(regWriteEnable_EXMEM_MEMWB),
		.instruction_EXMEM_MEMWB(instruction_EXMEM_MEMWB),
		.PC_EXMEM_MEMWB(PC_EXMEM_MEMWB),
		.regData2_EXMEM_out(regData2_EXMEM_out),
		.memType_EXMEM_out(memType_EXMEM_out),
		.memRead_EXMEM_MEMWB(memRead_EXMEM_MEMWB),
		.memWrite_EXMEM_out(memWrite_EXMEM_out),
		.execute_result_EXMEM_MEMWB(execute_result_EXMEM_MEMWB), 
		.ECALL_EXMEM_MEMWB(ECALL_EXMEM_MEMWB)

    );



	memory iMemory(
		///// INPUTS  /////
		.clk(clk),
		.rst_n(rst_n),
		.execute_result_EXMEM_MEMWB(execute_result_EXMEM_MEMWB),
		.memWrite_EXMEM_out(memWrite_EXMEM_out),
		.memRead_EXMEM_MEMWB(memRead_EXMEM_MEMWB),
		.regData2_EXMEM_out(regData2_EXMEM_out),
		.memType_EXMEM_out(memType_EXMEM_out),

		///// OUTPUTS  /////
		.memReadRst_MEMWB_in(memReadRst_MEMWB_in)
	
	);

	MEMWBpipelineReg iMEMWB_pipeline_reg(
		///// INPUTS  /////
		.clk(clk),
		.rst_n(rst_n),
		
		.stall_disable(1'b0),
		.flush(1'b0),

		///// PIPELINE INPUTS  /////
		.regWriteEnable_EXMEM_MEMWB(regWriteEnable_EXMEM_MEMWB),
		.instruction_EXMEM_MEMWB(instruction_EXMEM_MEMWB),
		.PC_EXMEM_MEMWB(PC_EXMEM_MEMWB),
		.execute_result_EXMEM_MEMWB(execute_result_EXMEM_MEMWB),
		.memRead_EXMEM_MEMWB(memRead_EXMEM_MEMWB),
		.memReadRst_MEMWB_in(memReadRst_MEMWB_in),
		.ECALL_EXMEM_MEMWB(ECALL_EXMEM_MEMWB),

		///// PIPELINE OUTPUTS  /////
		.regWriteEnable_MEMWB_out(regWriteEnable_MEMWB_out),
		.instruction_MEMWB_out(instruction_MEMWB_out),
		.PC_MEMWB_out(PC_MEMWB_out),
		.execute_result_MEMWB_out(execute_result_MEMWB_out),
		.memRead_MEMWB_out(memRead_MEMWB_out),
		.memReadRst_MEMWB_out(memReadRst_MEMWB_out),
		.ECALL_MEMWB_out(ECALL_MEMWB_out)

	);


	wb iWB(
        ///// INPUTS  /////
        .memReadRst_MEMWB_out(memReadRst_MEMWB_out),
        .memRead_MEMWB_out(memRead_MEMWB_out),
        .execute_result_MEMWB_out(execute_result_MEMWB_out),

        ///// OUTPUTS  /////
        .writeBackData(writeBackData)

        );

endmodule

`default_nettype wire
