module IM(clk,addr,rd_en,instr);

input clk;
input [15:0] addr;
input rd_en;			// asserted when instruction read desired

output reg [15:0] instr;	//output of insturction memory

reg [15:0]instr_mem[0:16383];

////////////////////////
// Instruction Memory //
////////////////////////
always @(negedge clk)
  if(rd_en) 
    instr <= instr_mem[addr];

/////////////////////////////
// Load Instruction Memory //
/////////////////////////////
initial begin
  $readmemh("HelloWorld.hex",instr_mem);
end

endmodule
