/*
    CS/ECE 552 Spring '23
    Eric Dubberstein, Joash Shankar

    LRU 256 input mux
*/
`default_nettype none
module LRUmux(
    // input
    index, stored_bits,
    
    // outputs
    data_out
    );

    input wire [7:0] index;
    output reg data_out;
    input wire [255:0] stored_bits;
	
	always@(*) begin
		case(index)
			8'd0: data_out = stored_bits[0];
			8'd1: data_out = stored_bits[1];
			8'd2: data_out = stored_bits[2];
			8'd3: data_out = stored_bits[3];
			8'd4: data_out = stored_bits[4];
			8'd5: data_out = stored_bits[5];
			8'd6: data_out = stored_bits[6];
			8'd7: data_out = stored_bits[7];
			8'd8: data_out = stored_bits[8];
			8'd9: data_out = stored_bits[9];
			8'd10: data_out = stored_bits[10];
			8'd11: data_out = stored_bits[11];
			8'd12: data_out = stored_bits[12];
			8'd13: data_out = stored_bits[13];
			8'd14: data_out = stored_bits[14];
			8'd15: data_out = stored_bits[15];
			8'd16: data_out = stored_bits[16];
			8'd17: data_out = stored_bits[17];
			8'd18: data_out = stored_bits[18];
			8'd19: data_out = stored_bits[19];
			8'd20: data_out = stored_bits[20];
			8'd21: data_out = stored_bits[21];
			8'd22: data_out = stored_bits[22];
			8'd23: data_out = stored_bits[23];
			8'd24: data_out = stored_bits[24];
			8'd25: data_out = stored_bits[25];
			8'd26: data_out = stored_bits[26];
			8'd27: data_out = stored_bits[27];
			8'd28: data_out = stored_bits[28];
			8'd29: data_out = stored_bits[29];
			8'd30: data_out = stored_bits[30];
			8'd31: data_out = stored_bits[31];
			8'd32: data_out = stored_bits[32];
			8'd33: data_out = stored_bits[33];
			8'd34: data_out = stored_bits[34];
			8'd35: data_out = stored_bits[35];
			8'd36: data_out = stored_bits[36];
			8'd37: data_out = stored_bits[37];
			8'd38: data_out = stored_bits[38];
			8'd39: data_out = stored_bits[39];
			8'd40: data_out = stored_bits[40];
			8'd41: data_out = stored_bits[41];
			8'd42: data_out = stored_bits[42];
			8'd43: data_out = stored_bits[43];
			8'd44: data_out = stored_bits[44];
			8'd45: data_out = stored_bits[45];
			8'd46: data_out = stored_bits[46];
			8'd47: data_out = stored_bits[47];
			8'd48: data_out = stored_bits[48];
			8'd49: data_out = stored_bits[49];
			8'd50: data_out = stored_bits[50];
			8'd51: data_out = stored_bits[51];
			8'd52: data_out = stored_bits[52];
			8'd53: data_out = stored_bits[53];
			8'd54: data_out = stored_bits[54];
			8'd55: data_out = stored_bits[55];
			8'd56: data_out = stored_bits[56];
			8'd57: data_out = stored_bits[57];
			8'd58: data_out = stored_bits[58];
			8'd59: data_out = stored_bits[59];
			8'd60: data_out = stored_bits[60];
			8'd61: data_out = stored_bits[61];
			8'd62: data_out = stored_bits[62];
			8'd63: data_out = stored_bits[63];
			8'd64: data_out = stored_bits[64];
			8'd65: data_out = stored_bits[65];
			8'd66: data_out = stored_bits[66];
			8'd67: data_out = stored_bits[67];
			8'd68: data_out = stored_bits[68];
			8'd69: data_out = stored_bits[69];
			8'd70: data_out = stored_bits[70];
			8'd71: data_out = stored_bits[71];
			8'd72: data_out = stored_bits[72];
			8'd73: data_out = stored_bits[73];
			8'd74: data_out = stored_bits[74];
			8'd75: data_out = stored_bits[75];
			8'd76: data_out = stored_bits[76];
			8'd77: data_out = stored_bits[77];
			8'd78: data_out = stored_bits[78];
			8'd79: data_out = stored_bits[79];
			8'd80: data_out = stored_bits[80];
			8'd81: data_out = stored_bits[81];
			8'd82: data_out = stored_bits[82];
			8'd83: data_out = stored_bits[83];
			8'd84: data_out = stored_bits[84];
			8'd85: data_out = stored_bits[85];
			8'd86: data_out = stored_bits[86];
			8'd87: data_out = stored_bits[87];
			8'd88: data_out = stored_bits[88];
			8'd89: data_out = stored_bits[89];
			8'd90: data_out = stored_bits[90];
			8'd91: data_out = stored_bits[91];
			8'd92: data_out = stored_bits[92];
			8'd93: data_out = stored_bits[93];
			8'd94: data_out = stored_bits[94];
			8'd95: data_out = stored_bits[95];
			8'd96: data_out = stored_bits[96];
			8'd97: data_out = stored_bits[97];
			8'd98: data_out = stored_bits[98];
			8'd99: data_out = stored_bits[99];
			8'd100: data_out = stored_bits[100];
			8'd101: data_out = stored_bits[101];
			8'd102: data_out = stored_bits[102];
			8'd103: data_out = stored_bits[103];
			8'd104: data_out = stored_bits[104];
			8'd105: data_out = stored_bits[105];
			8'd106: data_out = stored_bits[106];
			8'd107: data_out = stored_bits[107];
			8'd108: data_out = stored_bits[108];
			8'd109: data_out = stored_bits[109];
			8'd110: data_out = stored_bits[110];
			8'd111: data_out = stored_bits[111];
			8'd112: data_out = stored_bits[112];
			8'd113: data_out = stored_bits[113];
			8'd114: data_out = stored_bits[114];
			8'd115: data_out = stored_bits[115];
			8'd116: data_out = stored_bits[116];
			8'd117: data_out = stored_bits[117];
			8'd118: data_out = stored_bits[118];
			8'd119: data_out = stored_bits[119];
			8'd120: data_out = stored_bits[120];
			8'd121: data_out = stored_bits[121];
			8'd122: data_out = stored_bits[122];
			8'd123: data_out = stored_bits[123];
			8'd124: data_out = stored_bits[124];
			8'd125: data_out = stored_bits[125];
			8'd126: data_out = stored_bits[126];
			8'd127: data_out = stored_bits[127];
			8'd128: data_out = stored_bits[128];
			8'd129: data_out = stored_bits[129];
			8'd130: data_out = stored_bits[130];
			8'd131: data_out = stored_bits[131];
			8'd132: data_out = stored_bits[132];
			8'd133: data_out = stored_bits[133];
			8'd134: data_out = stored_bits[134];
			8'd135: data_out = stored_bits[135];
			8'd136: data_out = stored_bits[136];
			8'd137: data_out = stored_bits[137];
			8'd138: data_out = stored_bits[138];
			8'd139: data_out = stored_bits[139];
			8'd140: data_out = stored_bits[140];
			8'd141: data_out = stored_bits[141];
			8'd142: data_out = stored_bits[142];
			8'd143: data_out = stored_bits[143];
			8'd144: data_out = stored_bits[144];
			8'd145: data_out = stored_bits[145];
			8'd146: data_out = stored_bits[146];
			8'd147: data_out = stored_bits[147];
			8'd148: data_out = stored_bits[148];
			8'd149: data_out = stored_bits[149];
			8'd150: data_out = stored_bits[150];
			8'd151: data_out = stored_bits[151];
			8'd152: data_out = stored_bits[152];
			8'd153: data_out = stored_bits[153];
			8'd154: data_out = stored_bits[154];
			8'd155: data_out = stored_bits[155];
			8'd156: data_out = stored_bits[156];
			8'd157: data_out = stored_bits[157];
			8'd158: data_out = stored_bits[158];
			8'd159: data_out = stored_bits[159];
			8'd160: data_out = stored_bits[160];
			8'd161: data_out = stored_bits[161];
			8'd162: data_out = stored_bits[162];
			8'd163: data_out = stored_bits[163];
			8'd164: data_out = stored_bits[164];
			8'd165: data_out = stored_bits[165];
			8'd166: data_out = stored_bits[166];
			8'd167: data_out = stored_bits[167];
			8'd168: data_out = stored_bits[168];
			8'd169: data_out = stored_bits[169];
			8'd170: data_out = stored_bits[170];
			8'd171: data_out = stored_bits[171];
			8'd172: data_out = stored_bits[172];
			8'd173: data_out = stored_bits[173];
			8'd174: data_out = stored_bits[174];
			8'd175: data_out = stored_bits[175];
			8'd176: data_out = stored_bits[176];
			8'd177: data_out = stored_bits[177];
			8'd178: data_out = stored_bits[178];
			8'd179: data_out = stored_bits[179];
			8'd180: data_out = stored_bits[180];
			8'd181: data_out = stored_bits[181];
			8'd182: data_out = stored_bits[182];
			8'd183: data_out = stored_bits[183];
			8'd184: data_out = stored_bits[184];
			8'd185: data_out = stored_bits[185];
			8'd186: data_out = stored_bits[186];
			8'd187: data_out = stored_bits[187];
			8'd188: data_out = stored_bits[188];
			8'd189: data_out = stored_bits[189];
			8'd190: data_out = stored_bits[190];
			8'd191: data_out = stored_bits[191];
			8'd192: data_out = stored_bits[192];
			8'd193: data_out = stored_bits[193];
			8'd194: data_out = stored_bits[194];
			8'd195: data_out = stored_bits[195];
			8'd196: data_out = stored_bits[196];
			8'd197: data_out = stored_bits[197];
			8'd198: data_out = stored_bits[198];
			8'd199: data_out = stored_bits[199];
			8'd200: data_out = stored_bits[200];
			8'd201: data_out = stored_bits[201];
			8'd202: data_out = stored_bits[202];
			8'd203: data_out = stored_bits[203];
			8'd204: data_out = stored_bits[204];
			8'd205: data_out = stored_bits[205];
			8'd206: data_out = stored_bits[206];
			8'd207: data_out = stored_bits[207];
			8'd208: data_out = stored_bits[208];
			8'd209: data_out = stored_bits[209];
			8'd210: data_out = stored_bits[210];
			8'd211: data_out = stored_bits[211];
			8'd212: data_out = stored_bits[212];
			8'd213: data_out = stored_bits[213];
			8'd214: data_out = stored_bits[214];
			8'd215: data_out = stored_bits[215];
			8'd216: data_out = stored_bits[216];
			8'd217: data_out = stored_bits[217];
			8'd218: data_out = stored_bits[218];
			8'd219: data_out = stored_bits[219];
			8'd220: data_out = stored_bits[220];
			8'd221: data_out = stored_bits[221];
			8'd222: data_out = stored_bits[222];
			8'd223: data_out = stored_bits[223];
			8'd224: data_out = stored_bits[224];
			8'd225: data_out = stored_bits[225];
			8'd226: data_out = stored_bits[226];
			8'd227: data_out = stored_bits[227];
			8'd228: data_out = stored_bits[228];
			8'd229: data_out = stored_bits[229];
			8'd230: data_out = stored_bits[230];
			8'd231: data_out = stored_bits[231];
			8'd232: data_out = stored_bits[232];
			8'd233: data_out = stored_bits[233];
			8'd234: data_out = stored_bits[234];
			8'd235: data_out = stored_bits[235];
			8'd236: data_out = stored_bits[236];
			8'd237: data_out = stored_bits[237];
			8'd238: data_out = stored_bits[238];
			8'd239: data_out = stored_bits[239];
			8'd240: data_out = stored_bits[240];
			8'd241: data_out = stored_bits[241];
			8'd242: data_out = stored_bits[242];
			8'd243: data_out = stored_bits[243];
			8'd244: data_out = stored_bits[244];
			8'd245: data_out = stored_bits[245];
			8'd246: data_out = stored_bits[246];
			8'd247: data_out = stored_bits[247];
			8'd248: data_out = stored_bits[248];
			8'd249: data_out = stored_bits[249];
			8'd250: data_out = stored_bits[250];
			8'd251: data_out = stored_bits[251];
			8'd252: data_out = stored_bits[252];
			8'd253: data_out = stored_bits[253];
			8'd254: data_out = stored_bits[254];
			8'd255: data_out = stored_bits[255];
		endcase
	end

endmodule
`default_nettype wire
