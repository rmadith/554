module ALU(
    input [31:0] A, B,
    input [3:0] ALU_op,
    output out
);






endmodule
